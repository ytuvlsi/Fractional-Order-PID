magic
tech sky130A
magscale 1 2
timestamp 1729086831
<< nwell >>
rect 2954 1808 3544 2010
<< viali >>
rect 1730 3366 4202 3402
rect 1730 2434 1918 2468
rect 1608 1740 3412 1774
rect 3940 1580 3976 1866
rect 3736 -640 3776 -50
<< metal1 >>
rect 1716 3402 4214 3408
rect 1716 3366 1730 3402
rect 4202 3366 4214 3402
rect 1716 3360 4214 3366
rect 1716 3218 1752 3360
rect 4058 3308 4068 3328
rect 1790 3258 4068 3308
rect 1716 3200 1762 3218
rect 1728 2474 1762 3200
rect 1856 2586 1906 3258
rect 4058 3248 4068 3258
rect 4154 3248 4164 3328
rect 3044 2626 3054 2762
rect 3152 2626 3162 2762
rect 3288 2624 3298 2760
rect 3396 2624 3406 2760
rect 3522 2630 3532 2766
rect 3630 2630 3640 2766
rect 3758 2636 3768 2772
rect 3866 2636 3876 2772
rect 3990 2642 4000 2778
rect 4098 2642 4108 2778
rect 1800 2584 1906 2586
rect 1800 2520 1872 2584
rect 1862 2504 1872 2520
rect 1954 2504 1964 2584
rect 1718 2468 1930 2474
rect 1718 2434 1730 2468
rect 1918 2434 1930 2468
rect 1718 2428 1930 2434
rect 1728 2384 1762 2428
rect 1728 2382 2218 2384
rect 1610 2380 2218 2382
rect 1608 2312 2218 2380
rect 1608 2238 2120 2312
rect 2216 2238 2226 2312
rect 2382 2240 2392 2320
rect 2478 2240 2488 2320
rect 2616 2242 2626 2322
rect 2712 2242 2722 2322
rect 3166 2294 3176 2440
rect 3270 2294 3280 2440
rect 3406 2300 3416 2446
rect 3510 2300 3520 2446
rect 3640 2300 3650 2446
rect 3744 2300 3754 2446
rect 3878 2300 3888 2446
rect 3982 2300 3992 2446
rect 4114 2298 4124 2444
rect 4218 2298 4228 2444
rect 1608 2184 2218 2238
rect 1608 2182 1782 2184
rect 1608 1780 1712 2182
rect 1758 1900 1870 2100
rect 1952 1900 1962 2100
rect 2278 2034 2288 2124
rect 2360 2034 2370 2124
rect 2510 2038 2520 2128
rect 2592 2038 2602 2128
rect 2748 2042 2758 2132
rect 2830 2042 2840 2132
rect 3110 2100 3120 2180
rect 3198 2126 4072 2180
rect 3198 2100 3208 2126
rect 4062 2100 4072 2126
rect 4158 2100 4168 2180
rect 2000 1900 2170 1980
rect 2252 1978 2262 1980
rect 2252 1920 2692 1978
rect 2252 1900 2262 1920
rect 2682 1898 2692 1920
rect 2770 1898 2780 1978
rect 3602 1942 3802 1944
rect 1596 1774 3424 1780
rect 1596 1740 1608 1774
rect 3412 1740 3424 1774
rect 3590 1742 3600 1942
rect 3800 1878 3810 1942
rect 3800 1866 4052 1878
rect 3800 1744 3940 1866
rect 3800 1742 3810 1744
rect 1596 1734 3424 1740
rect 1160 1680 1360 1682
rect 1160 1632 2328 1680
rect 2678 1632 3860 1680
rect 1160 1078 1360 1632
rect 1710 1092 1720 1268
rect 1804 1092 1814 1268
rect 1950 1090 1960 1266
rect 2044 1090 2054 1266
rect 2190 1094 2200 1270
rect 2284 1094 2294 1270
rect 1158 878 1360 1078
rect 1160 350 1360 878
rect 2338 778 2684 960
rect 1602 600 1612 758
rect 1674 600 1684 758
rect 1840 598 1850 756
rect 1912 598 1922 756
rect 2076 602 2086 760
rect 2148 602 2158 760
rect 2328 600 2338 778
rect 2684 600 2694 778
rect 2870 606 2880 764
rect 2942 606 2952 764
rect 3102 608 3112 766
rect 3174 608 3184 766
rect 3338 608 3348 766
rect 3410 608 3420 766
rect 1946 384 1956 490
rect 2050 384 2060 490
rect 2338 402 2684 600
rect 3660 354 3860 1632
rect 3934 1580 3940 1744
rect 3976 1786 4052 1866
rect 4094 1818 4704 1866
rect 3976 1580 4096 1786
rect 3934 1568 3982 1580
rect 4142 1562 4152 1718
rect 4230 1562 4240 1718
rect 4382 1562 4392 1718
rect 4470 1562 4480 1718
rect 4016 790 4026 1014
rect 4110 790 4120 1014
rect 4260 780 4270 1004
rect 4354 780 4364 1004
rect 4620 804 4704 1818
rect 4792 1560 4802 1758
rect 5002 1560 5012 1758
rect 4800 1558 5000 1560
rect 4620 556 4658 804
rect 4082 438 4092 556
rect 4408 464 4658 556
rect 4914 464 4924 804
rect 4408 460 4708 464
rect 4408 438 4418 460
rect 1160 298 2328 350
rect 2694 302 3862 354
rect 3660 298 3860 302
rect 3414 6 3424 86
rect 3622 56 3632 86
rect 3622 6 4362 56
rect 3422 4 4362 6
rect 3422 -16 3622 4
rect 3892 -2 4362 4
rect 3472 -56 3576 -16
rect 3892 -20 4098 -2
rect 3730 -50 3782 -38
rect 3730 -54 3736 -50
rect 3348 -408 3358 -254
rect 3450 -408 3460 -254
rect 3492 -680 3548 -56
rect 3626 -252 3736 -54
rect 3776 -54 3782 -50
rect 3776 -252 3894 -54
rect 3936 -190 3946 -62
rect 4038 -190 4048 -62
rect 3596 -406 3606 -252
rect 3610 -408 3620 -406
rect 3902 -254 3912 -252
rect 3626 -636 3736 -408
rect 3730 -640 3736 -636
rect 3776 -418 3830 -408
rect 3906 -418 3916 -254
rect 4066 -416 4076 -252
rect 4152 -416 4162 -252
rect 3776 -636 3894 -418
rect 3776 -640 3782 -636
rect 3730 -652 3782 -640
rect 4280 -680 4362 -2
rect 3420 -702 3620 -680
rect 3880 -702 4362 -680
rect 3420 -756 4362 -702
<< via1 >>
rect 4068 3248 4154 3328
rect 3054 2626 3152 2762
rect 3298 2624 3396 2760
rect 3532 2630 3630 2766
rect 3768 2636 3866 2772
rect 4000 2642 4098 2778
rect 1872 2504 1954 2584
rect 2120 2238 2216 2312
rect 2392 2240 2478 2320
rect 2626 2242 2712 2322
rect 3176 2294 3270 2440
rect 3416 2300 3510 2446
rect 3650 2300 3744 2446
rect 3888 2300 3982 2446
rect 4124 2298 4218 2444
rect 1870 1900 1952 2100
rect 2288 2034 2360 2124
rect 2520 2038 2592 2128
rect 2758 2042 2830 2132
rect 3120 2100 3198 2180
rect 4072 2100 4158 2180
rect 2170 1900 2252 1980
rect 2692 1898 2770 1978
rect 3600 1742 3800 1942
rect 1720 1092 1804 1268
rect 1960 1090 2044 1266
rect 2200 1094 2284 1270
rect 1612 600 1674 758
rect 1850 598 1912 756
rect 2086 602 2148 760
rect 2338 600 2684 778
rect 2880 606 2942 764
rect 3112 608 3174 766
rect 3348 608 3410 766
rect 1956 384 2050 490
rect 4152 1562 4230 1718
rect 4392 1562 4470 1718
rect 4026 790 4110 1014
rect 4270 780 4354 1004
rect 4802 1560 5002 1758
rect 4092 438 4408 556
rect 4658 464 4914 804
rect 3424 6 3622 86
rect 3358 -408 3450 -254
rect 3946 -190 4038 -62
rect 3606 -406 3736 -252
rect 3620 -408 3736 -406
rect 3736 -408 3776 -252
rect 3776 -254 3902 -252
rect 3776 -408 3906 -254
rect 3830 -418 3906 -408
rect 4076 -416 4152 -252
<< metal2 >>
rect 4068 3328 4340 3338
rect 4154 3248 4340 3328
rect 4068 3240 4340 3248
rect 4068 3238 4154 3240
rect 2126 2778 4104 2788
rect 2126 2772 4000 2778
rect 2126 2766 3768 2772
rect 2126 2762 3532 2766
rect 2126 2626 3054 2762
rect 3152 2760 3532 2762
rect 3152 2626 3298 2760
rect 2126 2624 3298 2626
rect 3396 2630 3532 2760
rect 3630 2636 3768 2766
rect 3866 2642 4000 2772
rect 4098 2642 4104 2778
rect 3866 2636 4104 2642
rect 3630 2630 4104 2636
rect 3396 2624 4104 2630
rect 2126 2620 4104 2624
rect 1872 2592 1954 2594
rect 1870 2584 1954 2592
rect 1870 2504 1872 2584
rect 1870 2494 1954 2504
rect 1870 2100 1952 2494
rect 2126 2322 2322 2620
rect 3054 2616 3152 2620
rect 3298 2614 3396 2620
rect 3416 2450 3510 2456
rect 3650 2450 3744 2456
rect 3888 2450 3982 2456
rect 4124 2450 4218 2454
rect 3166 2446 4218 2450
rect 3166 2440 3416 2446
rect 2392 2322 2478 2330
rect 2626 2322 2712 2332
rect 2120 2320 2626 2322
rect 2120 2312 2392 2320
rect 2216 2240 2392 2312
rect 2478 2242 2626 2320
rect 3166 2294 3176 2440
rect 3270 2300 3416 2440
rect 3510 2300 3650 2446
rect 3744 2300 3888 2446
rect 3982 2444 4218 2446
rect 3982 2300 4124 2444
rect 3270 2298 4124 2300
rect 3270 2294 4218 2298
rect 3166 2290 4218 2294
rect 3176 2284 3270 2290
rect 2478 2240 2712 2242
rect 2216 2238 2322 2240
rect 2120 2236 2322 2238
rect 2120 2228 2216 2236
rect 2392 2230 2478 2240
rect 2626 2232 2712 2240
rect 3120 2180 3200 2190
rect 2758 2138 2830 2142
rect 2288 2132 2832 2138
rect 2288 2128 2758 2132
rect 2288 2124 2520 2128
rect 2360 2038 2520 2124
rect 2592 2042 2758 2128
rect 2830 2042 2832 2132
rect 3198 2100 3200 2180
rect 3120 2090 3200 2100
rect 2592 2038 2832 2042
rect 2360 2034 2832 2038
rect 2288 2022 2832 2034
rect 2170 1980 2252 1990
rect 1952 1900 2170 1980
rect 1870 1890 1952 1900
rect 2170 1890 2252 1900
rect 1720 1272 1804 1278
rect 1960 1272 2044 1276
rect 2200 1272 2284 1280
rect 1720 1270 2292 1272
rect 1720 1268 2200 1270
rect 1804 1266 2200 1268
rect 1804 1092 1960 1266
rect 1720 1090 1960 1092
rect 2044 1094 2200 1266
rect 2284 1094 2292 1270
rect 2044 1090 2292 1094
rect 1720 1086 2292 1090
rect 1720 1082 1804 1086
rect 1960 1080 2044 1086
rect 2200 1084 2284 1086
rect 2442 788 2576 2022
rect 2692 1980 2770 1988
rect 3122 1980 3200 2090
rect 2692 1978 3200 1980
rect 2770 1898 3200 1978
rect 3600 1942 3800 1952
rect 2692 1888 2770 1898
rect 3600 1732 3800 1742
rect 3856 1720 4008 2290
rect 4124 2288 4218 2290
rect 4072 2180 4158 2190
rect 4262 2180 4340 3240
rect 4158 2100 4342 2180
rect 4072 2088 4342 2100
rect 4802 1766 5002 1768
rect 4800 1758 5002 1766
rect 4800 1756 4802 1758
rect 4152 1720 4230 1728
rect 3856 1718 4230 1720
rect 4392 1718 4470 1728
rect 3856 1562 4152 1718
rect 4230 1562 4392 1718
rect 4470 1564 4800 1718
rect 4470 1562 4802 1564
rect 3856 1560 4802 1562
rect 5002 1560 5004 1718
rect 4152 1558 4470 1560
rect 4152 1552 4230 1558
rect 4392 1552 4470 1558
rect 4800 1554 5002 1560
rect 4802 1550 5002 1554
rect 4026 1014 4110 1024
rect 4020 790 4026 1012
rect 4270 1012 4354 1014
rect 4110 1004 4360 1012
rect 4110 790 4270 1004
rect 2338 778 2684 788
rect 1612 766 1674 768
rect 2086 766 2148 770
rect 1612 760 2338 766
rect 1612 758 2086 760
rect 1674 756 2086 758
rect 1674 600 1850 756
rect 1612 598 1850 600
rect 1912 602 2086 756
rect 2148 602 2338 760
rect 1912 600 2338 602
rect 4020 780 4270 790
rect 4354 780 4360 1004
rect 2880 766 2942 774
rect 3112 766 3174 776
rect 3348 766 3410 776
rect 4020 772 4360 780
rect 4658 804 4914 814
rect 4270 770 4354 772
rect 2684 764 3112 766
rect 2684 606 2880 764
rect 2942 608 3112 764
rect 3174 608 3348 766
rect 3410 608 3414 766
rect 2942 606 3414 608
rect 2684 600 3414 606
rect 1912 598 3414 600
rect 1612 596 3414 598
rect 1612 590 1674 596
rect 1850 588 1912 596
rect 2086 592 2148 596
rect 2338 590 2684 596
rect 4092 556 4408 566
rect 1956 498 2050 500
rect 1944 490 2056 498
rect 1944 384 1956 490
rect 2050 384 2056 490
rect 1944 96 2056 384
rect 3946 438 4092 556
rect 4658 454 4914 464
rect 3946 428 4408 438
rect 1944 86 3622 96
rect 1944 6 3424 86
rect 1944 -4 3622 6
rect 3946 -62 4102 428
rect 4038 -190 4102 -62
rect 3946 -200 4038 -190
rect 3606 -244 3902 -242
rect 3358 -250 3450 -244
rect 3606 -250 3906 -244
rect 3356 -252 3906 -250
rect 4076 -252 4152 -242
rect 3356 -254 3606 -252
rect 3902 -254 4076 -252
rect 3356 -408 3358 -254
rect 3450 -406 3606 -254
rect 3450 -408 3620 -406
rect 3358 -418 3450 -408
rect 3606 -416 3830 -408
rect 3620 -418 3830 -416
rect 3906 -416 4076 -254
rect 3906 -418 4152 -416
rect 3830 -422 4152 -418
rect 3830 -428 3906 -422
rect 4076 -426 4152 -422
<< via2 >>
rect 3600 1742 3800 1942
rect 4800 1564 4802 1756
rect 4802 1564 4998 1756
rect 4658 464 4914 804
<< metal3 >>
rect 3590 1944 3810 1947
rect 3590 1942 3836 1944
rect 3590 1742 3600 1942
rect 3800 1742 3836 1942
rect 3590 1737 3836 1742
rect 3620 -252 3836 1737
rect 4790 1756 5008 1761
rect 4790 1564 4800 1756
rect 4998 1564 5008 1756
rect 4790 1559 5008 1564
rect 4648 804 4924 809
rect 4648 464 4658 804
rect 4914 464 4924 804
rect 4648 459 4924 464
rect 3610 -408 3620 -252
rect 3902 -408 3912 -252
<< via3 >>
rect 4800 1564 4998 1756
rect 4658 464 4914 804
rect 3620 -408 3902 -252
<< metal4 >>
rect 5536 4106 6184 4108
rect 4806 3878 6186 4106
rect 4806 1757 5014 3878
rect 5536 3494 6184 3878
rect 4799 1756 5014 1757
rect 4799 1564 4800 1756
rect 4998 1564 5014 1756
rect 4799 1563 5014 1564
rect 4806 1554 5014 1563
rect 4657 804 4915 805
rect 4657 794 4658 804
rect 4656 466 4658 794
rect 4657 464 4658 466
rect 4914 794 4915 804
rect 4914 466 5254 794
rect 4914 464 4915 466
rect 4657 463 4915 464
rect 3619 -252 3903 -251
rect 3619 -408 3620 -252
rect 3902 -408 3903 -252
rect 3619 -409 3903 -408
use sky130_fd_pr__cap_mim_m3_1_XFFB5V  XC2
timestamp 1729082712
transform -1 0 6452 0 -1 1444
box -1286 -2240 1286 2240
use sky130_fd_pr__pfet_01v8_F6U8HA  XM1
timestamp 1729082712
transform 1 0 1824 0 1 2917
box -226 -519 226 519
use sky130_fd_pr__pfet_01v8_FEZMTC  XM2
timestamp 1729082712
transform 1 0 2494 0 1 2617
box -462 -819 462 819
use sky130_fd_pr__pfet_01v8_FGZ9KC  XM3
timestamp 1729082712
transform 1 0 1999 0 1 991
box -521 -819 521 819
use sky130_fd_pr__pfet_01v8_FGZ9KC  XM4
timestamp 1729082712
transform 1 0 3023 0 1 991
box -521 -819 521 819
use sky130_fd_pr__nfet_01v8_92UYLD  XM5
timestamp 1729082712
transform 1 0 3523 0 1 -350
box -285 -510 285 510
use sky130_fd_pr__nfet_01v8_92UYLD  XM6
timestamp 1729082712
transform 1 0 3987 0 1 -350
box -285 -510 285 510
use sky130_fd_pr__pfet_01v8_NQ9489  XM7
timestamp 1729082712
transform 1 0 3636 0 1 2719
box -698 -719 698 719
use sky130_fd_pr__nfet_01v8_BGD4RZ  XM8
timestamp 1729082712
transform 1 0 4248 0 1 1186
box -344 -810 344 810
<< labels >>
flabel metal1 1728 2184 1928 2384 0 FreeSans 256 0 0 0 VDD
port 3 nsew
flabel metal1 1758 1900 1958 2100 0 FreeSans 256 0 0 0 IBIAS
port 5 nsew
flabel metal1 1158 878 1358 1078 0 FreeSans 256 0 0 0 VN
port 0 nsew
flabel metal1 3660 880 3860 1080 0 FreeSans 256 0 0 0 VP
port 1 nsew
flabel metal1 3602 1744 3802 1944 0 FreeSans 256 0 0 0 GND
port 2 nsew
flabel metal1 4800 1558 5000 1758 0 FreeSans 256 0 0 0 VOUT
port 4 nsew
<< end >>
