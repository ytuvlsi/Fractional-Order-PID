magic
tech sky130A
magscale 1 2
timestamp 1729011116
<< viali >>
rect 6330 3150 6530 3184
rect 5948 806 5984 1058
rect 6864 802 6900 1054
rect 40 -126 78 202
rect 5950 -300 5986 -48
rect 6864 -302 6900 -50
rect 8584 -1024 8784 -970
rect 4112 -1532 4148 -1172
<< metal1 >>
rect 6330 3190 6530 3562
rect 5374 3189 6542 3190
rect 5330 3188 6542 3189
rect 7432 3189 7482 3190
rect 7432 3188 7524 3189
rect 5330 3184 7524 3188
rect 5330 3150 6330 3184
rect 6530 3150 7524 3184
rect 5330 3142 7524 3150
rect 5330 3140 5422 3142
rect 6330 3140 7524 3142
rect 5330 3002 5376 3140
rect 5330 2958 5378 3002
rect 5600 2598 5660 3044
rect 5810 3042 5896 3088
rect 6060 2598 6120 3052
rect 6210 3032 6220 3094
rect 6280 3032 6290 3094
rect 6330 3002 6530 3140
rect 6578 3028 6588 3104
rect 6658 3028 6668 3104
rect 5600 2518 6120 2598
rect 5600 2112 5660 2518
rect 6060 2372 6120 2518
rect 6290 2112 6566 3002
rect 6740 2112 6800 3052
rect 6954 3042 7040 3088
rect 7200 2112 7260 3052
rect 7478 3008 7524 3140
rect 7476 2960 7524 3008
rect 5600 1958 5660 2004
rect 5812 1998 5822 2064
rect 5890 1998 5900 2064
rect 6326 2004 6526 2112
rect 6290 2000 6564 2004
rect 5812 1914 5898 1960
rect 6740 1958 6800 2004
rect 6956 1990 6966 2056
rect 7030 1990 7040 2056
rect 6954 1914 7040 1960
rect 7200 1958 7260 2004
rect 7710 1806 7720 2004
rect 7854 1806 7998 2004
rect 7798 1804 7998 1806
rect 596 1600 5818 1644
rect 7030 1600 7454 1648
rect 7538 1640 12256 1648
rect 7458 1600 12256 1640
rect 172 534 372 610
rect 510 578 520 656
rect 602 578 612 656
rect 1030 536 1114 1600
rect 1560 1476 1570 1560
rect 1662 1476 1672 1560
rect 2058 536 2142 1600
rect 2628 596 2638 674
rect 2720 596 2730 674
rect 3198 536 3282 1600
rect 3684 1480 3694 1560
rect 3778 1480 3788 1560
rect 4226 536 4310 1600
rect 4744 572 4754 650
rect 4836 572 4846 650
rect 5406 536 5490 1600
rect 5806 1496 5816 1562
rect 5890 1496 5900 1562
rect 6956 1488 6966 1554
rect 7030 1488 7040 1554
rect 5942 1058 5990 1070
rect 5942 806 5948 1058
rect 5984 980 5990 1058
rect 6858 1054 6906 1066
rect 6858 1036 6864 1054
rect 5984 900 6442 980
rect 5984 806 5990 900
rect 5942 794 5990 806
rect 172 486 632 534
rect 832 488 5820 536
rect 172 410 372 486
rect 3830 238 3840 266
rect 34 202 84 214
rect 34 134 40 202
rect -2 128 40 134
rect 78 128 84 202
rect 150 200 3840 238
rect 4002 238 4012 266
rect 4002 200 4592 238
rect 150 192 4592 200
rect 4828 196 5122 488
rect 150 148 196 192
rect -22 -64 -12 128
rect 80 -64 90 128
rect -2 -126 40 -64
rect 78 -126 84 -64
rect -2 -138 84 -126
rect -2 -1156 66 -138
rect 114 -798 124 -700
rect 224 -798 234 -700
rect 318 -888 384 192
rect 468 52 478 152
rect 582 52 592 152
rect 670 -898 736 192
rect 868 138 914 192
rect 828 -800 838 -702
rect 938 -800 948 -702
rect 1028 -896 1094 192
rect 1188 30 1198 130
rect 1302 30 1312 130
rect 1394 -896 1460 192
rect 1582 140 1628 192
rect 1542 -800 1552 -702
rect 1652 -800 1662 -702
rect 1768 -894 1834 192
rect 1892 26 1902 126
rect 2006 26 2016 126
rect 2106 -898 2172 192
rect 2300 140 2346 192
rect 2260 -800 2270 -702
rect 2370 -800 2380 -702
rect 2474 -898 2540 192
rect 2622 30 2632 130
rect 2736 30 2746 130
rect 2810 -898 2876 192
rect 3014 142 3060 192
rect 2976 -800 2986 -702
rect 3086 -800 3096 -702
rect 3168 -902 3234 192
rect 3332 34 3342 134
rect 3446 34 3456 134
rect 3526 -902 3592 192
rect 3730 152 3776 192
rect 3690 -800 3700 -702
rect 3800 -800 3810 -702
rect 3902 -896 3968 192
rect 4052 28 4062 128
rect 4166 28 4176 128
rect 4242 -904 4308 192
rect 4446 164 4592 192
rect 4446 -166 4818 164
rect 4446 -518 4752 -166
rect 4860 -518 4870 -166
rect 4446 -728 4818 -518
rect 4408 -814 4418 -728
rect 4506 -814 4818 -728
rect 4446 -840 4818 -814
rect 5298 -900 5382 228
rect 5872 120 5920 612
rect 5944 -48 5992 -36
rect 5944 -300 5950 -48
rect 5986 -66 5992 -48
rect 5986 -288 5988 -66
rect 6070 -288 6080 -66
rect 6348 -130 6442 900
rect 6776 814 6786 1036
rect 6858 802 6864 814
rect 6900 802 6906 1054
rect 6858 790 6906 802
rect 6932 112 6980 604
rect 7458 536 7542 1600
rect 8004 570 8014 638
rect 8094 570 8104 638
rect 8596 536 8680 1600
rect 9062 1488 9072 1566
rect 9156 1488 9166 1566
rect 9572 536 9656 1600
rect 10120 582 10130 650
rect 10210 582 10220 650
rect 10710 536 10794 1600
rect 11176 1482 11186 1560
rect 11270 1482 11280 1560
rect 11686 536 11770 1600
rect 12238 578 12248 646
rect 12328 578 12338 646
rect 7030 524 12066 536
rect 12486 534 12686 594
rect 7030 502 12004 524
rect 7030 488 11940 502
rect 12230 492 12686 534
rect 6858 -50 6906 -38
rect 6858 -124 6864 -50
rect 6796 -130 6864 -124
rect 6348 -210 6864 -130
rect 5986 -300 5992 -288
rect 5944 -312 5992 -300
rect 6796 -302 6864 -210
rect 6900 -302 6906 -50
rect 6796 -314 6906 -302
rect 6796 -670 6896 -314
rect 6790 -774 6800 -670
rect 6886 -774 6896 -670
rect 7486 -898 7570 236
rect 7728 196 8022 488
rect 12486 394 12686 492
rect 8834 246 8844 268
rect 8420 202 8844 246
rect 9006 246 9016 268
rect 9006 202 12650 246
rect 8420 200 12650 202
rect 8028 120 8412 164
rect 8028 -50 8274 120
rect 8418 -50 8428 120
rect 8028 -320 8412 -50
rect 7998 -760 8008 -320
rect 8100 -760 8412 -320
rect 8028 -838 8412 -760
rect 8532 -902 8598 200
rect 8672 -830 8682 -666
rect 8806 -830 8816 -666
rect 8896 -902 8962 200
rect 9030 -60 9040 110
rect 9184 -60 9194 110
rect 9254 -898 9320 200
rect 9386 -824 9396 -660
rect 9520 -824 9530 -660
rect 9624 -898 9690 200
rect 9742 -60 9752 110
rect 9896 -60 9906 110
rect 9958 -910 10024 200
rect 10108 -820 10118 -656
rect 10242 -820 10252 -656
rect 10326 -906 10392 200
rect 10454 -62 10464 108
rect 10608 -62 10618 108
rect 10682 -906 10748 200
rect 10820 -818 10830 -654
rect 10954 -818 10964 -654
rect 11020 -902 11086 200
rect 11168 -62 11178 108
rect 11322 -62 11332 108
rect 11406 -906 11472 200
rect 11536 -818 11546 -654
rect 11670 -818 11680 -654
rect 11740 -910 11806 200
rect 11878 -60 11888 110
rect 12032 -60 12042 110
rect 12092 -902 12158 200
rect 12258 -820 12268 -656
rect 12392 -820 12402 -656
rect 12468 -902 12534 200
rect 12616 -62 12626 108
rect 12770 -62 12780 108
rect 8572 -970 8796 -964
rect 8572 -1024 8584 -970
rect 8784 -1024 8796 -970
rect 8572 -1030 8796 -1024
rect -2 -1172 4156 -1156
rect 4742 -1168 4804 -1166
rect 5482 -1168 5544 -1162
rect 5828 -1168 5890 -1166
rect 6054 -1168 6064 -1112
rect -2 -1400 4112 -1172
rect 0 -1442 4112 -1400
rect 1175 -1532 4112 -1442
rect 4148 -1246 4156 -1172
rect 4274 -1208 6064 -1168
rect 6720 -1168 6730 -1112
rect 6720 -1208 8508 -1168
rect 4274 -1218 8508 -1208
rect 4148 -1396 4268 -1246
rect 4148 -1532 4156 -1396
rect 1175 -1602 4156 -1532
rect 4146 -1606 4156 -1602
rect 4282 -1606 4292 -1396
rect 4372 -2278 4434 -1218
rect 4532 -2198 4542 -2026
rect 4652 -2198 4662 -2026
rect 4742 -2278 4804 -1218
rect 4892 -1600 4902 -1390
rect 5028 -1600 5038 -1390
rect 5090 -2278 5152 -1218
rect 5256 -2192 5266 -2020
rect 5376 -2192 5386 -2020
rect 5482 -2278 5544 -1218
rect 5612 -1602 5622 -1392
rect 5748 -1602 5758 -1392
rect 5828 -2278 5890 -1218
rect 5968 -2186 5978 -2014
rect 6088 -2186 6098 -2014
rect 6170 -2278 6232 -1218
rect 6324 -1602 6334 -1392
rect 6460 -1602 6470 -1392
rect 6528 -2278 6590 -1218
rect 6688 -2184 6698 -2012
rect 6808 -2184 6818 -2012
rect 6898 -2278 6960 -1218
rect 7036 -1602 7046 -1392
rect 7172 -1602 7182 -1392
rect 7234 -2278 7296 -1218
rect 7398 -2186 7408 -2014
rect 7518 -2186 7528 -2014
rect 7600 -2278 7662 -1218
rect 7754 -1604 7764 -1394
rect 7890 -1604 7900 -1394
rect 7968 -2278 8030 -1218
rect 8114 -2184 8124 -2012
rect 8234 -2184 8244 -2012
rect 8328 -2278 8390 -1218
rect 8468 -1604 8478 -1394
rect 8604 -1604 8614 -1394
rect 8940 -2200 8950 -1998
rect 9056 -2000 9066 -1998
rect 9056 -2200 9200 -2000
rect 4276 -2328 8508 -2278
rect 5090 -2330 5152 -2328
rect 6170 -2334 6232 -2328
rect 6528 -2334 6590 -2328
rect 6898 -2330 6960 -2328
rect 7234 -2334 7296 -2328
rect 7600 -2334 7662 -2328
rect 7968 -2332 8030 -2328
rect 8328 -2330 8390 -2328
<< via1 >>
rect 6220 3032 6280 3094
rect 6588 3028 6658 3104
rect 5822 1998 5890 2064
rect 6966 1990 7030 2056
rect 7720 1806 7854 2004
rect 520 578 602 656
rect 1570 1476 1662 1560
rect 2638 596 2720 674
rect 3694 1480 3778 1560
rect 4754 572 4836 650
rect 5816 1496 5890 1562
rect 6966 1488 7030 1554
rect 3840 200 4002 266
rect -12 -64 40 128
rect 40 -64 78 128
rect 78 -64 80 128
rect 124 -798 224 -700
rect 478 52 582 152
rect 838 -800 938 -702
rect 1198 30 1302 130
rect 1552 -800 1652 -702
rect 1902 26 2006 126
rect 2270 -800 2370 -702
rect 2632 30 2736 130
rect 2986 -800 3086 -702
rect 3342 34 3446 134
rect 3700 -800 3800 -702
rect 4062 28 4166 128
rect 4752 -518 4860 -166
rect 4418 -814 4506 -728
rect 5988 -288 6070 -66
rect 6786 814 6864 1036
rect 6864 814 6868 1036
rect 8014 570 8094 638
rect 9072 1488 9156 1566
rect 10130 582 10210 650
rect 11186 1482 11270 1560
rect 12248 578 12328 646
rect 6800 -774 6886 -670
rect 8844 202 9006 268
rect 8274 -50 8418 120
rect 8008 -760 8100 -320
rect 8682 -830 8806 -666
rect 9040 -60 9184 110
rect 9396 -824 9520 -660
rect 9752 -60 9896 110
rect 10118 -820 10242 -656
rect 10464 -62 10608 108
rect 10830 -818 10954 -654
rect 11178 -62 11322 108
rect 11546 -818 11670 -654
rect 11888 -60 12032 110
rect 12268 -820 12392 -656
rect 12626 -62 12770 108
rect 8584 -1024 8784 -970
rect 6064 -1208 6720 -1112
rect 4156 -1606 4282 -1396
rect 4542 -2198 4652 -2026
rect 4902 -1600 5028 -1390
rect 5266 -2192 5376 -2020
rect 5622 -1602 5748 -1392
rect 5978 -2186 6088 -2014
rect 6334 -1602 6460 -1392
rect 6698 -2184 6808 -2012
rect 7046 -1602 7172 -1392
rect 7408 -2186 7518 -2014
rect 7764 -1604 7890 -1394
rect 8124 -2184 8234 -2012
rect 8478 -1604 8604 -1394
rect 8950 -2200 9056 -1998
<< metal2 >>
rect 6588 3108 6658 3114
rect 6220 3104 6660 3108
rect 6220 3094 6588 3104
rect 6280 3032 6588 3094
rect 6220 3028 6588 3032
rect 6658 3028 6660 3104
rect 6220 3020 6660 3028
rect 6588 3018 6658 3020
rect 5822 2064 5890 2074
rect 5816 1998 5822 2000
rect 6966 2056 7030 2066
rect 5890 1998 5894 2000
rect 5816 1570 5894 1998
rect 7720 2004 7854 2014
rect 7030 1990 7720 1996
rect 6966 1806 7720 1990
rect 7854 1806 7858 1996
rect 6966 1802 7858 1806
rect 6966 1572 7030 1802
rect 7720 1796 7854 1802
rect 9072 1572 9156 1576
rect 1570 1562 5898 1570
rect 1570 1560 5816 1562
rect 1662 1480 3694 1560
rect 3778 1496 5816 1560
rect 5890 1496 5898 1562
rect 3778 1480 5898 1496
rect 1662 1476 5898 1480
rect 6954 1566 11270 1572
rect 6954 1554 9072 1566
rect 6954 1488 6966 1554
rect 7030 1488 9072 1554
rect 9156 1560 11270 1566
rect 9156 1488 11186 1560
rect 6954 1482 11186 1488
rect 6954 1476 11270 1482
rect 1570 1462 5898 1476
rect 11186 1472 11270 1476
rect 6786 1036 6868 1046
rect 6236 814 6786 890
rect 6236 804 6868 814
rect 6236 796 6812 804
rect 2638 674 2720 684
rect 520 660 602 666
rect 520 656 2638 660
rect 602 596 2638 656
rect 2720 650 4838 660
rect 2720 596 4754 650
rect 602 578 4754 596
rect 520 572 4754 578
rect 4836 572 4838 650
rect 520 568 4838 572
rect 3840 266 4002 276
rect 3840 190 4002 200
rect 478 152 582 162
rect -10 138 478 140
rect -12 128 478 138
rect 80 52 478 128
rect 3342 140 3446 144
rect 582 138 4164 140
rect 582 134 4166 138
rect 582 130 3342 134
rect 582 52 1198 130
rect 80 30 1198 52
rect 1302 126 2632 130
rect 1302 30 1902 126
rect 80 26 618 30
rect 1198 20 1302 30
rect 2006 30 2632 126
rect 2736 34 3342 130
rect 3446 128 4166 134
rect 3446 34 4062 128
rect 2736 30 4062 34
rect 1902 16 2006 26
rect 2632 20 2736 30
rect 3342 24 3446 30
rect 4062 18 4166 28
rect -12 -74 80 -64
rect 4364 -580 4490 568
rect 4754 562 4836 568
rect 5988 -58 6070 -56
rect 6236 -58 6332 796
rect 7450 660 7622 664
rect 7450 658 8050 660
rect 10130 658 10210 660
rect 7450 650 12330 658
rect 7450 638 10130 650
rect 7450 570 8014 638
rect 8094 582 10130 638
rect 10210 646 12330 650
rect 10210 582 12248 646
rect 8094 578 12248 582
rect 12328 578 12330 646
rect 8094 570 12330 578
rect 7450 562 12330 570
rect 7450 560 8094 562
rect 7450 552 8050 560
rect 7450 -58 7622 552
rect 8844 268 9006 278
rect 8844 192 9006 202
rect 8274 128 8418 130
rect 4750 -66 7622 -58
rect 4750 -166 5988 -66
rect 4750 -378 4752 -166
rect 4860 -288 5988 -166
rect 6070 -288 7622 -66
rect 8264 120 12774 128
rect 8264 -50 8274 120
rect 8418 110 12774 120
rect 8418 -50 9040 110
rect 8264 -60 9040 -50
rect 9184 -60 9752 110
rect 9896 108 11888 110
rect 9896 -60 10464 108
rect 8264 -62 10464 -60
rect 10608 -62 11178 108
rect 11322 -60 11888 108
rect 12032 108 12774 110
rect 12032 -60 12626 108
rect 11322 -62 12626 -60
rect 12770 -62 12774 108
rect 8264 -70 12774 -62
rect 10464 -72 10608 -70
rect 11178 -72 11322 -70
rect 12626 -72 12770 -70
rect 4860 -378 7622 -288
rect 8008 -320 8100 -310
rect 4752 -528 4860 -518
rect 4364 -670 6904 -580
rect 4364 -682 6800 -670
rect 124 -700 224 -690
rect 116 -798 124 -714
rect 838 -702 938 -692
rect 224 -798 838 -714
rect 116 -800 838 -798
rect 1552 -702 1652 -692
rect 938 -800 1552 -714
rect 2270 -702 2370 -692
rect 1652 -800 2270 -714
rect 2986 -702 3086 -692
rect 2370 -800 2986 -714
rect 3700 -702 3800 -692
rect 3086 -800 3700 -714
rect 3800 -718 4452 -714
rect 3800 -728 4506 -718
rect 3800 -800 4418 -728
rect 124 -808 224 -800
rect 838 -810 938 -800
rect 1552 -810 1652 -800
rect 2270 -810 2370 -800
rect 2986 -810 3086 -800
rect 3700 -810 3800 -800
rect 6886 -760 8008 -670
rect 8544 -654 12394 -644
rect 8544 -656 10830 -654
rect 8544 -660 10118 -656
rect 8544 -666 9396 -660
rect 8100 -760 8108 -670
rect 6886 -772 8108 -760
rect 6800 -784 6886 -774
rect 4418 -824 4506 -814
rect 8544 -830 8682 -666
rect 8806 -824 9396 -666
rect 9520 -820 10118 -660
rect 10242 -818 10830 -656
rect 10954 -818 11546 -654
rect 11670 -656 12394 -654
rect 11670 -818 12268 -656
rect 10242 -820 12268 -818
rect 12392 -820 12394 -656
rect 9520 -824 12394 -820
rect 8806 -830 12394 -824
rect 8544 -844 12394 -830
rect 8544 -970 8822 -844
rect 8544 -1024 8584 -970
rect 8784 -1024 8822 -970
rect 6064 -1112 6720 -1102
rect 6064 -1218 6720 -1208
rect 4902 -1382 5028 -1380
rect 8544 -1382 8822 -1024
rect 4154 -1390 8822 -1382
rect 4154 -1396 4902 -1390
rect 4154 -1606 4156 -1396
rect 4282 -1600 4902 -1396
rect 5028 -1392 8822 -1390
rect 5028 -1600 5622 -1392
rect 4282 -1602 5622 -1600
rect 5748 -1602 6334 -1392
rect 6460 -1602 7046 -1392
rect 7172 -1394 8822 -1392
rect 7172 -1602 7764 -1394
rect 4282 -1604 7764 -1602
rect 7890 -1604 8478 -1394
rect 8604 -1604 8822 -1394
rect 4282 -1606 8822 -1604
rect 4154 -1618 8822 -1606
rect 8950 -1994 9056 -1988
rect 8114 -1996 9062 -1994
rect 4542 -1998 9062 -1996
rect 4542 -2012 8950 -1998
rect 4542 -2014 6698 -2012
rect 4542 -2020 5978 -2014
rect 4542 -2026 5266 -2020
rect 4652 -2192 5266 -2026
rect 5376 -2186 5978 -2020
rect 6088 -2184 6698 -2014
rect 6808 -2014 8124 -2012
rect 6808 -2184 7408 -2014
rect 6088 -2186 7408 -2184
rect 7518 -2184 8124 -2014
rect 8234 -2184 8950 -2012
rect 7518 -2186 8950 -2184
rect 5376 -2192 8950 -2186
rect 4652 -2198 8950 -2192
rect 4542 -2200 8950 -2198
rect 9056 -2200 9062 -1998
rect 4542 -2208 9062 -2200
rect 4542 -2210 8234 -2208
rect 8950 -2210 9056 -2208
<< via2 >>
rect 3840 200 4002 266
rect 8844 202 9006 268
rect 6064 -1208 6720 -1112
<< metal3 >>
rect 3830 268 4012 271
rect 6064 268 6722 270
rect 8834 268 9016 273
rect 3830 266 8844 268
rect 3830 200 3840 266
rect 4002 202 8844 266
rect 9006 202 9016 268
rect 4002 200 9016 202
rect 3830 195 4012 200
rect 6064 -1107 6722 200
rect 8834 197 9016 200
rect 6054 -1112 6730 -1107
rect 6054 -1208 6064 -1112
rect 6720 -1208 6730 -1112
rect 6054 -1213 6730 -1208
use sky130_fd_pr__nfet_01v8_T5X68Y  XMb1
timestamp 1728988403
transform 1 0 6387 0 1 -1748
box -2315 -710 2315 710
use sky130_fd_pr__nfet_01v8_T5X68Y  XMb2
timestamp 1728988403
transform 1 0 2321 0 1 -338
box -2315 -710 2315 710
use sky130_fd_pr__nfet_01v8_T5X68Y  XMb3
timestamp 1728988403
transform 1 0 10523 0 1 -340
box -2315 -710 2315 710
use sky130_fd_pr__nfet_01v8_6NWCSU  XMn1
timestamp 1728988403
transform 1 0 3206 0 1 1064
box -2812 -710 2812 710
use sky130_fd_pr__nfet_01v8_2Z49SJ  XMn2
timestamp 1728988403
transform 1 0 7530 0 1 -338
box -696 -710 696 710
use sky130_fd_pr__nfet_01v8_2Z49SJ  XMn3
timestamp 1728988403
transform 1 0 5322 0 1 -338
box -696 -710 696 710
use sky130_fd_pr__nfet_01v8_6NWCSU  XMn4
timestamp 1728988403
transform 1 0 9638 0 1 1065
box -2812 -710 2812 710
use sky130_fd_pr__pfet_01v8_UQS8UX  XMp1
timestamp 1728988403
transform 1 0 5855 0 1 2501
box -625 -719 625 719
use sky130_fd_pr__pfet_01v8_UQS8UX  XMp2
timestamp 1728988403
transform 1 0 6999 0 1 2501
box -625 -719 625 719
<< labels >>
flabel metal1 6330 3362 6530 3562 0 FreeSans 256 0 0 0 VDD
port 1 nsew
flabel metal1 172 410 372 610 0 FreeSans 256 0 0 0 VP
port 5 nsew
flabel metal1 12486 394 12686 594 0 FreeSans 256 0 0 0 VN
port 4 nsew
flabel metal1 -2 -1400 198 -1200 0 FreeSans 256 0 0 0 VSS
port 3 nsew
flabel metal1 9000 -2200 9200 -2000 0 FreeSans 256 0 0 0 IBIAS
port 0 nsew
flabel metal1 7798 1804 7998 2004 0 FreeSans 256 0 0 0 IOUT
port 2 nsew
<< end >>
