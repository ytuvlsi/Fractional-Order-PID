magic
tech sky130A
magscale 1 2
timestamp 1729526722
<< metal1 >>
rect 5796 14006 76218 14010
rect 88076 14006 88812 14010
rect 5796 12730 5998 14006
rect 7262 14000 88812 14006
rect 7262 12750 80024 14000
rect 81810 12750 88812 14000
rect 7262 12730 88812 12750
rect 5796 12728 76218 12730
rect 85152 12226 85162 12440
rect 86104 12226 86114 12440
rect 12284 11216 12294 11418
rect 12498 11216 12508 11418
rect 25262 11216 25272 11414
rect 25476 11216 25486 11414
rect 38236 11178 38246 11382
rect 38468 11178 38478 11382
rect 51224 11138 51234 11344
rect 51438 11138 51448 11344
rect 64150 11064 64160 11266
rect 64352 11064 64362 11266
rect 77102 11024 77112 11228
rect 77326 11024 77336 11228
rect 68726 10708 69000 10716
rect 55796 10686 56000 10702
rect 29824 10670 30044 10678
rect 16856 10648 17082 10654
rect 16856 10302 16948 10648
rect 17594 10302 17604 10648
rect 29824 10340 29954 10670
rect 30598 10340 30608 10670
rect 3200 10202 4188 10206
rect 3200 9804 4746 10202
rect 3200 612 4188 9804
rect 16856 9802 17082 10302
rect 17488 9808 17498 10044
rect 17730 9808 17740 10044
rect 29824 9804 30044 10340
rect 42814 10294 42894 10624
rect 43614 10294 43624 10624
rect 55796 10304 55866 10686
rect 56600 10304 56610 10686
rect 68726 10306 68800 10708
rect 69416 10306 69426 10708
rect 30486 9780 30496 9986
rect 30700 9780 30710 9986
rect 42814 9768 43022 10294
rect 43470 9744 43480 9956
rect 43686 9744 43696 9956
rect 55796 9726 56000 10304
rect 56414 9870 56614 9872
rect 56402 9670 56412 9870
rect 56616 9670 56626 9870
rect 68726 9652 69000 10306
rect 69350 9630 69360 9838
rect 69564 9630 69574 9838
rect 82032 9828 82334 9832
rect 81674 9610 82334 9828
rect 4328 7580 4338 8256
rect 5724 7580 5734 8256
rect 17894 7596 17904 8250
rect 20042 7596 20052 8250
rect 30896 7560 30906 8214
rect 33044 7560 33054 8214
rect 43848 7514 43858 8168
rect 45996 7514 46006 8168
rect 56846 7442 56856 8096
rect 58994 7442 59004 8096
rect 69858 7414 69868 8068
rect 72006 7414 72016 8068
rect 4944 6432 4954 6914
rect 5320 6432 5330 6914
rect 13370 6908 27802 6912
rect 39416 6908 39680 6914
rect 52428 6908 52642 6914
rect 5988 6886 7798 6888
rect 13370 6886 56656 6908
rect 5974 6832 56656 6886
rect 65326 6832 65602 6834
rect 5974 6804 70600 6832
rect 5974 6796 81804 6804
rect 5974 6498 79990 6796
rect 5988 6202 7798 6498
rect 13370 6478 79990 6498
rect 27800 6474 79990 6478
rect 56168 6398 79990 6474
rect 70580 6388 79990 6398
rect 81798 6388 81808 6796
rect 70580 6372 81804 6388
rect 5978 5592 5988 6202
rect 7794 5592 7804 6202
rect 12270 5062 12280 5262
rect 12480 5062 12490 5262
rect 25204 5062 25214 5262
rect 25414 5062 25424 5262
rect 38176 5002 38186 5202
rect 38386 5002 38396 5202
rect 51144 4948 51154 5154
rect 51358 4948 51368 5154
rect 64116 4930 64126 5134
rect 64310 4930 64320 5134
rect 77068 4946 77078 5150
rect 77292 4946 77302 5150
rect 78592 4952 78602 5400
rect 79600 4952 79610 5400
rect 4514 3662 4524 3866
rect 4770 3662 4780 3866
rect 16784 3652 16794 3854
rect 17038 3652 17048 3854
rect 17458 3666 17468 3868
rect 17706 3666 17716 3868
rect 29726 3650 29736 3858
rect 29992 3650 30002 3858
rect 30408 3608 30418 3816
rect 30646 3608 30656 3816
rect 42680 3594 42690 3800
rect 42936 3594 42946 3800
rect 43412 3550 43422 3760
rect 43670 3550 43680 3760
rect 55686 3536 55696 3738
rect 55940 3536 55950 3738
rect 56382 3534 56392 3742
rect 56624 3534 56634 3742
rect 68646 3520 68656 3722
rect 68908 3520 68918 3722
rect 69318 3550 69328 3756
rect 69580 3550 69590 3756
rect 81612 3536 81622 3738
rect 81850 3536 81860 3738
rect 4860 820 4870 2100
rect 8002 820 8012 2100
rect 13350 1054 13550 1254
rect 17902 820 17912 2100
rect 21044 820 21054 2100
rect 26302 1056 26502 1256
rect 30900 762 30910 2042
rect 34042 762 34052 2042
rect 39248 998 39448 1198
rect 43864 720 43874 2000
rect 47006 720 47016 2000
rect 52252 946 52452 1146
rect 56842 782 56852 1974
rect 60004 782 60014 1974
rect 65222 922 65422 1122
rect 69860 806 69870 1998
rect 73022 806 73032 1998
rect 78160 940 78360 1140
rect 3200 608 16800 612
rect 82032 608 82334 9610
rect 82790 8604 82800 9986
rect 83598 8604 83608 9986
rect 88076 5996 88812 12730
rect 87004 4800 88794 4808
rect 86554 4698 88794 4800
rect 86522 4524 86532 4698
rect 86782 4596 88794 4698
rect 86782 4524 86792 4596
rect 87004 3400 88794 4596
rect 86812 808 86822 2210
rect 87800 808 87810 2210
rect 3200 -450 83514 608
rect 85132 -96 85142 142
rect 85634 -96 85644 142
rect 3200 -466 29548 -450
rect 3200 -1010 16792 -466
rect 17202 -1002 29548 -466
rect 17202 -1010 17212 -1002
rect 29538 -1006 29548 -1002
rect 30024 -456 83514 -450
rect 30024 -462 85786 -456
rect 30024 -468 81622 -462
rect 30024 -472 68530 -468
rect 30024 -1002 42526 -472
rect 30024 -1006 30034 -1002
rect 42516 -1004 42526 -1002
rect 42988 -474 68530 -472
rect 42988 -1002 55516 -474
rect 42988 -1004 42998 -1002
rect 55506 -1004 55516 -1002
rect 55968 -1000 68530 -474
rect 68930 -1000 81622 -468
rect 82004 -1000 85786 -462
rect 55968 -1002 82016 -1000
rect 55968 -1004 55978 -1002
rect 81964 -1006 82016 -1002
rect 3200 -1014 16800 -1010
rect 85776 -1014 85786 -1000
rect 86262 -1014 86272 -456
rect 69252 -1200 69262 -1186
rect 4400 -1202 69262 -1200
rect 4400 -1204 30332 -1202
rect 4400 -1786 4532 -1204
rect 4394 -1804 4532 -1786
rect 4874 -1206 30332 -1204
rect 4874 -1804 17392 -1206
rect 4394 -1814 17392 -1804
rect 17848 -1798 30332 -1206
rect 30832 -1204 69262 -1202
rect 30832 -1206 56320 -1204
rect 30832 -1798 43352 -1206
rect 17848 -1810 43352 -1798
rect 43806 -1806 56320 -1206
rect 56798 -1806 69262 -1204
rect 69728 -1806 69738 -1186
rect 43806 -1810 69736 -1806
rect 17848 -1814 69736 -1810
rect 4394 -2404 69736 -1814
<< via1 >>
rect 5998 12730 7262 14006
rect 80024 12750 81810 14000
rect 85162 12226 86104 12440
rect 12294 11216 12498 11418
rect 25272 11216 25476 11414
rect 38246 11178 38468 11382
rect 51234 11138 51438 11344
rect 64160 11064 64352 11266
rect 77112 11024 77326 11228
rect 16948 10302 17594 10648
rect 29954 10340 30598 10670
rect 17498 9808 17730 10044
rect 42894 10294 43614 10624
rect 55866 10304 56600 10686
rect 68800 10306 69416 10708
rect 30496 9780 30700 9986
rect 43480 9744 43686 9956
rect 56412 9670 56616 9870
rect 69360 9630 69564 9838
rect 4338 7580 5724 8256
rect 17904 7596 20042 8250
rect 30906 7560 33044 8214
rect 43858 7514 45996 8168
rect 56856 7442 58994 8096
rect 69868 7414 72006 8068
rect 4954 6432 5320 6914
rect 79990 6388 81798 6796
rect 5988 5592 7794 6202
rect 12280 5062 12480 5262
rect 25214 5062 25414 5262
rect 38186 5002 38386 5202
rect 51154 4948 51358 5154
rect 64126 4930 64310 5134
rect 77078 4946 77292 5150
rect 78602 4952 79600 5400
rect 4524 3662 4770 3866
rect 16794 3652 17038 3854
rect 17468 3666 17706 3868
rect 29736 3650 29992 3858
rect 30418 3608 30646 3816
rect 42690 3594 42936 3800
rect 43422 3550 43670 3760
rect 55696 3536 55940 3738
rect 56392 3534 56624 3742
rect 68656 3520 68908 3722
rect 69328 3550 69580 3756
rect 81622 3536 81850 3738
rect 4870 820 8002 2100
rect 17912 820 21044 2100
rect 30910 762 34042 2042
rect 43874 720 47006 2000
rect 56852 782 60004 1974
rect 69870 806 73022 1998
rect 82800 8604 83598 9986
rect 86532 4524 86782 4698
rect 86822 808 87800 2210
rect 85142 -96 85634 142
rect 16792 -1010 17202 -466
rect 29548 -1006 30024 -450
rect 42526 -1004 42988 -472
rect 55516 -1004 55968 -474
rect 68530 -1000 68930 -468
rect 81622 -1000 82004 -462
rect 85786 -1014 86262 -456
rect 4532 -1804 4874 -1204
rect 17392 -1814 17848 -1206
rect 30332 -1798 30832 -1202
rect 43352 -1810 43806 -1206
rect 56320 -1806 56798 -1204
rect 69262 -1806 69728 -1186
<< metal2 >>
rect 5998 14006 7262 14016
rect 80024 14000 81810 14010
rect 80024 12740 81810 12750
rect 5998 12720 7262 12730
rect 85162 12440 86104 12450
rect 85162 12216 86104 12226
rect 12294 11418 12498 11428
rect 12294 11206 12498 11216
rect 25272 11414 25476 11424
rect 25272 11206 25476 11216
rect 38246 11382 38468 11392
rect 38246 11168 38468 11178
rect 51234 11344 51438 11354
rect 51234 11128 51438 11138
rect 64160 11266 64352 11276
rect 64160 11054 64352 11064
rect 77112 11228 77326 11238
rect 77112 11014 77326 11024
rect 68800 10708 69416 10718
rect 55866 10686 56600 10696
rect 29954 10670 30598 10680
rect 16948 10648 17594 10658
rect 29954 10330 30598 10340
rect 42894 10624 43614 10634
rect 16948 10292 17594 10302
rect 55866 10294 56600 10304
rect 68800 10296 69416 10306
rect 42894 10284 43614 10294
rect 17498 10044 17730 10054
rect 17498 9798 17730 9808
rect 30496 9986 30700 9996
rect 82800 9986 83598 9996
rect 30496 9770 30700 9780
rect 43480 9956 43686 9966
rect 43480 9734 43686 9744
rect 56412 9870 56616 9880
rect 56412 9660 56616 9670
rect 69360 9838 69564 9848
rect 69360 9620 69564 9630
rect 82800 8594 83598 8604
rect 4338 8256 5724 8266
rect 17904 8250 20042 8260
rect 17904 7586 20042 7596
rect 30906 8214 33044 8224
rect 4338 7570 5724 7580
rect 30906 7550 33044 7560
rect 43858 8168 45996 8178
rect 43858 7504 45996 7514
rect 56856 8096 58994 8106
rect 56856 7432 58994 7442
rect 69868 8068 72006 8078
rect 4954 6914 5320 6924
rect 13280 6914 13434 7418
rect 26150 6914 26394 7414
rect 69868 7404 72006 7414
rect 39152 6914 39384 7382
rect 52104 6914 52370 7346
rect 64974 6914 65308 7268
rect 77944 6916 78242 7228
rect 65342 6914 65590 6916
rect 77430 6914 78280 6916
rect 4948 6432 4954 6914
rect 5320 6912 26470 6914
rect 26648 6912 78280 6914
rect 5320 6432 78280 6912
rect 4948 6428 78280 6432
rect 4954 6422 5320 6428
rect 77430 6218 78280 6428
rect 79982 6796 81798 6808
rect 79982 6388 79990 6796
rect 79982 6372 81798 6388
rect 5988 6202 7794 6212
rect 77430 5702 82756 6218
rect 5988 5582 7794 5592
rect 78602 5400 79600 5410
rect 12280 5262 12480 5272
rect 12280 5052 12480 5062
rect 25214 5262 25414 5272
rect 25214 5052 25414 5062
rect 38186 5202 38386 5212
rect 38186 4992 38386 5002
rect 51154 5154 51358 5164
rect 77078 5150 77292 5160
rect 51154 4938 51358 4948
rect 64126 5134 64310 5144
rect 77078 4936 77292 4946
rect 78602 4942 79600 4952
rect 64126 4920 64310 4930
rect 4524 3866 4770 3876
rect 17468 3868 17706 3878
rect 4770 3662 4772 3866
rect 4524 3652 4772 3662
rect 4654 -1194 4772 3652
rect 16794 3854 17038 3864
rect 17468 3656 17706 3666
rect 16794 3642 17038 3652
rect 4870 2100 8002 2110
rect 4870 810 8002 820
rect 16794 -456 16912 3642
rect 16792 -466 17202 -456
rect 16792 -1020 17202 -1010
rect 4532 -1204 4874 -1194
rect 17570 -1196 17706 3656
rect 29736 3858 29992 3868
rect 29736 3640 29992 3650
rect 30418 3816 30646 3826
rect 17912 2100 21044 2110
rect 17912 810 21044 820
rect 29740 -440 29874 3640
rect 30418 3598 30646 3608
rect 42690 3800 42936 3810
rect 29548 -450 30024 -440
rect 29548 -1016 30024 -1006
rect 30534 -1192 30644 3598
rect 42690 3584 42936 3594
rect 43422 3760 43670 3770
rect 30910 2042 34042 2052
rect 30910 752 34042 762
rect 42690 -462 42816 3584
rect 43670 3550 43672 3758
rect 69328 3756 69580 3766
rect 43422 3540 43672 3550
rect 42526 -472 42988 -462
rect 42526 -1014 42988 -1004
rect 4532 -1814 4874 -1804
rect 17392 -1206 17848 -1196
rect 30332 -1202 30832 -1192
rect 43530 -1196 43672 3540
rect 55696 3738 55940 3748
rect 55696 3526 55940 3536
rect 56392 3742 56624 3752
rect 43874 2000 47006 2010
rect 43874 710 47006 720
rect 55696 -464 55818 3526
rect 56392 3524 56624 3534
rect 55516 -474 55968 -464
rect 55516 -1014 55968 -1004
rect 56496 -1194 56624 3524
rect 68656 3722 68908 3732
rect 69328 3540 69580 3550
rect 81622 3738 81850 3748
rect 68656 3510 68908 3520
rect 56852 1974 60004 1984
rect 56852 772 60004 782
rect 68658 -458 68786 3510
rect 68530 -468 68930 -458
rect 68530 -1010 68930 -1000
rect 69452 -1176 69574 3540
rect 81622 3526 81850 3536
rect 69870 1998 73022 2008
rect 69870 796 73022 806
rect 81622 -452 81740 3526
rect 85142 142 85634 152
rect 85142 -106 85634 -96
rect 85786 -446 86102 12216
rect 86532 4698 86782 4708
rect 86532 4514 86782 4524
rect 86822 2210 87800 2220
rect 86822 798 87800 808
rect 81622 -462 82004 -452
rect 81622 -1010 82004 -1000
rect 85786 -456 86262 -446
rect 85786 -1024 86262 -1014
rect 69262 -1186 69728 -1176
rect 30332 -1808 30832 -1798
rect 43352 -1206 43806 -1196
rect 17392 -1824 17848 -1814
rect 43352 -1820 43806 -1810
rect 56320 -1204 56798 -1194
rect 56320 -1816 56798 -1806
rect 69262 -1816 69728 -1806
<< via2 >>
rect 5998 12730 7262 14006
rect 80024 12750 81810 14000
rect 12294 11216 12498 11418
rect 25272 11216 25476 11414
rect 38246 11178 38468 11382
rect 51234 11138 51438 11344
rect 64160 11064 64352 11266
rect 77112 11024 77326 11228
rect 16948 10302 17594 10648
rect 29954 10340 30598 10670
rect 42894 10294 43614 10624
rect 55866 10304 56600 10686
rect 68800 10306 69416 10708
rect 17498 9808 17730 10044
rect 30496 9780 30700 9986
rect 43480 9744 43686 9956
rect 56412 9670 56616 9870
rect 69360 9630 69564 9838
rect 82800 8604 83598 9986
rect 4338 7580 5724 8256
rect 17904 7596 20042 8250
rect 30906 7560 33044 8214
rect 43858 7514 45996 8168
rect 56856 7442 58994 8096
rect 69868 7414 72006 8068
rect 79990 6388 81798 6796
rect 5988 5592 7794 6202
rect 12280 5062 12480 5262
rect 25214 5062 25414 5262
rect 38186 5002 38386 5202
rect 51154 4948 51358 5154
rect 64126 4930 64310 5134
rect 77078 4946 77292 5150
rect 78602 4952 79600 5400
rect 4870 820 8002 2100
rect 17912 820 21044 2100
rect 30910 762 34042 2042
rect 43874 720 47006 2000
rect 56852 782 60004 1974
rect 69870 806 73022 1998
rect 85142 -96 85634 142
rect 86532 4524 86782 4698
rect 86822 808 87800 2210
<< metal3 >>
rect 5988 14006 7272 14011
rect 5988 12730 5998 14006
rect 7262 12730 7272 14006
rect 80014 14000 81820 14005
rect 80014 12750 80024 14000
rect 81810 12750 81820 14000
rect 80014 12745 81820 12750
rect 5988 12725 7272 12730
rect 85400 11800 86240 11802
rect 12294 11423 14602 11600
rect 12284 11418 14602 11423
rect 25272 11419 27604 11602
rect 12284 11216 12294 11418
rect 12498 11216 14602 11418
rect 25262 11414 27604 11419
rect 25262 11216 25272 11414
rect 25476 11216 27604 11414
rect 38246 11387 40602 11600
rect 12284 11211 12508 11216
rect 13598 10196 14600 11216
rect 25262 11211 25486 11216
rect 16938 10648 17604 10653
rect 16938 10302 16948 10648
rect 17594 10302 17604 10648
rect 16938 10297 17604 10302
rect 13598 10049 17732 10196
rect 26576 10190 27604 11216
rect 38236 11382 40602 11387
rect 38236 11178 38246 11382
rect 38468 11178 40602 11382
rect 51234 11596 53600 11602
rect 51234 11349 53606 11596
rect 51224 11344 53606 11349
rect 38236 11173 38478 11178
rect 29944 10670 30608 10675
rect 29944 10340 29954 10670
rect 30598 10340 30608 10670
rect 29944 10335 30608 10340
rect 13598 10044 17740 10049
rect 13598 9808 17498 10044
rect 17730 9808 17740 10044
rect 13598 9803 17740 9808
rect 26576 9991 30706 10190
rect 39596 10144 40600 11178
rect 51224 11138 51234 11344
rect 51438 11138 53606 11344
rect 64160 11271 66600 11406
rect 78602 11404 86240 11800
rect 78598 11402 86240 11404
rect 51224 11133 51448 11138
rect 42884 10624 43624 10629
rect 42884 10294 42894 10624
rect 43614 10294 43624 10624
rect 42884 10289 43624 10294
rect 52604 10196 53606 11138
rect 64150 11266 66600 11271
rect 64150 11064 64160 11266
rect 64352 11064 66600 11266
rect 77112 11233 86240 11402
rect 64150 11059 64362 11064
rect 55856 10686 56610 10691
rect 55856 10304 55866 10686
rect 56600 10304 56610 10686
rect 55856 10299 56610 10304
rect 26576 9986 30710 9991
rect 13598 9604 17732 9803
rect 26576 9780 30496 9986
rect 30700 9780 30710 9986
rect 26576 9775 30710 9780
rect 39596 9956 43734 10144
rect 4328 8256 5734 8261
rect 4328 7580 4338 8256
rect 5724 7580 5734 8256
rect 4328 7575 5734 7580
rect 4332 2105 5730 7575
rect 5978 6202 7804 6207
rect 5978 5592 5988 6202
rect 7794 5592 7804 6202
rect 5978 5587 7804 5592
rect 13598 5400 14600 9604
rect 26576 9600 30706 9775
rect 39596 9744 43480 9956
rect 43686 9744 43734 9956
rect 39596 9604 43734 9744
rect 52602 9870 56634 10196
rect 52602 9670 56412 9870
rect 56616 9670 56634 9870
rect 17894 8250 20052 8255
rect 17894 7596 17904 8250
rect 20042 7596 20052 8250
rect 17894 7591 20052 7596
rect 12280 5267 14602 5400
rect 12270 5262 14602 5267
rect 12270 5062 12280 5262
rect 12480 5062 14602 5262
rect 12270 5057 12490 5062
rect 17904 2105 20034 7591
rect 26576 5404 27604 9600
rect 30896 8214 33054 8219
rect 30896 7560 30906 8214
rect 33044 7560 33054 8214
rect 30896 7555 33054 7560
rect 25212 5267 27610 5404
rect 25204 5262 27610 5267
rect 25204 5062 25214 5262
rect 25414 5062 27610 5262
rect 25204 5057 25424 5062
rect 4332 2100 8012 2105
rect 4332 828 4870 2100
rect 4350 822 4870 828
rect 4860 820 4870 822
rect 8002 1788 8012 2100
rect 17902 2100 21054 2105
rect 17902 1788 17912 2100
rect 8002 822 17912 1788
rect 8002 820 8012 822
rect 4860 815 8012 820
rect 17902 820 17912 822
rect 21044 1788 21054 2100
rect 30906 2047 33036 7555
rect 39596 7444 40600 9604
rect 52602 9596 56634 9670
rect 65596 10142 66600 11064
rect 77102 11228 86240 11233
rect 77102 11024 77112 11228
rect 77326 11026 86240 11228
rect 77326 11024 79600 11026
rect 77102 11019 77336 11024
rect 68790 10708 69426 10713
rect 68790 10306 68800 10708
rect 69416 10306 69426 10708
rect 68790 10301 69426 10306
rect 65596 9838 69604 10142
rect 65596 9630 69360 9838
rect 69564 9630 69604 9838
rect 43848 8168 46006 8173
rect 43848 7514 43858 8168
rect 45996 7514 46006 8168
rect 43848 7509 46006 7514
rect 39594 6516 40600 7444
rect 39596 5400 40600 6516
rect 38186 5207 40600 5400
rect 38176 5202 40600 5207
rect 38176 5002 38186 5202
rect 38386 5002 40600 5202
rect 38176 4997 38396 5002
rect 30900 2042 34052 2047
rect 30900 1788 30910 2042
rect 21044 822 30910 1788
rect 21044 820 21054 822
rect 17902 815 21054 820
rect 17904 798 20034 815
rect 30900 762 30910 822
rect 34042 1788 34052 2042
rect 43876 2005 46006 7509
rect 52604 5404 53606 9596
rect 65596 9570 69604 9630
rect 56846 8096 59004 8101
rect 56846 7442 56856 8096
rect 58994 7442 59004 8096
rect 56846 7437 59004 7442
rect 51190 5159 53606 5404
rect 51144 5154 53606 5159
rect 51144 4948 51154 5154
rect 51358 4950 53606 5154
rect 51358 4948 51368 4950
rect 51144 4943 51368 4948
rect 43864 2000 47016 2005
rect 43864 1788 43874 2000
rect 34042 822 43874 1788
rect 34042 762 34052 822
rect 30900 757 34052 762
rect 30906 736 33036 757
rect 43864 720 43874 822
rect 47006 1788 47016 2000
rect 56856 1979 58986 7437
rect 65596 5392 66600 9570
rect 69858 8068 72016 8073
rect 69858 7414 69868 8068
rect 72006 7414 72016 8068
rect 69858 7409 72016 7414
rect 64144 5139 66600 5392
rect 64116 5134 66600 5139
rect 64116 4930 64126 5134
rect 64310 4930 66600 5134
rect 64116 4926 66600 4930
rect 64116 4925 64320 4926
rect 69870 2003 72000 7409
rect 78598 5405 79598 11024
rect 82790 9986 83608 9991
rect 82790 8604 82800 9986
rect 83598 8604 83608 9986
rect 82790 8599 83608 8604
rect 79980 6796 81808 6801
rect 79980 6388 79990 6796
rect 81798 6388 81808 6796
rect 79980 6383 81808 6388
rect 78592 5400 79610 5405
rect 78592 5392 78602 5400
rect 77078 5155 78602 5392
rect 77068 5150 78602 5155
rect 77068 4946 77078 5150
rect 77292 4952 78602 5150
rect 79600 4952 79610 5400
rect 77292 4948 79610 4952
rect 77292 4946 77302 4948
rect 78592 4947 79610 4948
rect 77068 4941 77302 4946
rect 69860 1998 73032 2003
rect 56842 1974 60014 1979
rect 56842 1788 56852 1974
rect 47006 822 56852 1788
rect 47006 720 47016 822
rect 56842 782 56852 822
rect 60004 1788 60014 1974
rect 69860 1788 69870 1998
rect 60004 822 69870 1788
rect 60004 782 60014 822
rect 69860 806 69870 822
rect 73022 1788 73032 1998
rect 82526 1788 82536 2194
rect 73022 822 82536 1788
rect 73022 806 73032 822
rect 69860 801 73032 806
rect 82526 792 82536 822
rect 83514 792 83524 2194
rect 56842 777 60014 782
rect 56856 756 58986 777
rect 43864 715 47016 720
rect 43876 696 46006 715
rect 85400 147 86240 11026
rect 86522 4698 86792 4703
rect 86522 4524 86532 4698
rect 86782 4524 86792 4698
rect 86522 4519 86792 4524
rect 86812 2210 87810 2215
rect 86812 808 86822 2210
rect 87800 808 87810 2210
rect 86812 803 87810 808
rect 85132 142 86240 147
rect 85132 -96 85142 142
rect 85634 -94 86240 142
rect 85634 -96 85644 -94
rect 85132 -101 85644 -96
<< via3 >>
rect 5998 12730 7262 14006
rect 80024 12750 81810 14000
rect 16948 10302 17594 10648
rect 29954 10340 30598 10670
rect 42894 10294 43614 10624
rect 55866 10304 56600 10686
rect 5988 5592 7794 6202
rect 68800 10306 69416 10708
rect 82800 8604 83598 9986
rect 79990 6388 81798 6796
rect 78602 4952 79600 5400
rect 82536 792 83514 2194
rect 86532 4524 86782 4698
rect 86822 808 87800 2210
<< metal4 >>
rect 5997 14006 7263 14007
rect 5997 13994 5998 14006
rect 5988 12730 5998 13994
rect 7262 12730 7263 14006
rect 5988 12729 7263 12730
rect 79990 14001 81800 14016
rect 79990 14000 81811 14001
rect 79990 12750 80024 14000
rect 81810 12750 81811 14000
rect 79990 12749 81811 12750
rect 5988 6203 7262 12729
rect 16858 10710 55860 10712
rect 16858 10708 69426 10710
rect 16858 10686 68800 10708
rect 16858 10670 55866 10686
rect 16858 10648 29954 10670
rect 16858 10302 16948 10648
rect 17594 10340 29954 10648
rect 30598 10624 55866 10670
rect 30598 10340 42894 10624
rect 17594 10302 42894 10340
rect 16858 10294 42894 10302
rect 43614 10304 55866 10624
rect 56600 10306 68800 10686
rect 69416 10306 69426 10708
rect 56600 10304 69426 10306
rect 43614 10294 69426 10304
rect 16858 9802 69426 10294
rect 55798 9728 69426 9802
rect 5987 6202 7795 6203
rect 5987 5592 5988 6202
rect 7794 5592 7795 6202
rect 5987 5591 7795 5592
rect 68798 5402 69412 9728
rect 79990 6797 81800 12749
rect 87120 9996 87794 10002
rect 82800 9987 87814 9996
rect 82799 9986 87814 9987
rect 82799 8604 82800 9986
rect 83598 8604 87814 9986
rect 82799 8603 83599 8604
rect 79989 6796 81800 6797
rect 79989 6388 79990 6796
rect 81798 6388 81800 6796
rect 79989 6387 81799 6388
rect 68798 5400 79604 5402
rect 68798 5000 78602 5400
rect 78601 4952 78602 5000
rect 79600 5398 79604 5400
rect 79600 4952 87004 5398
rect 78601 4951 79601 4952
rect 86532 4699 86780 4952
rect 86531 4698 86783 4699
rect 86531 4524 86532 4698
rect 86782 4524 86783 4698
rect 86531 4523 86783 4524
rect 87120 2211 87794 8604
rect 86821 2210 87801 2211
rect 86821 2198 86822 2210
rect 82536 2195 86822 2198
rect 82535 2194 86822 2195
rect 82535 792 82536 2194
rect 83514 808 86822 2194
rect 87800 2198 87801 2210
rect 87800 808 87802 2198
rect 83514 792 87802 808
rect 82535 791 83515 792
use ota3  X1
timestamp 1729011116
transform 1 0 4372 0 1 9412
box -22 -2458 12838 3562
use ota3  X2
timestamp 1729011116
transform 1 0 17338 0 1 9412
box -22 -2458 12838 3562
use ota3  X3
timestamp 1729011116
transform 1 0 30326 0 1 9374
box -22 -2458 12838 3562
use ota3  X4
timestamp 1729011116
transform 1 0 43312 0 1 9336
box -22 -2458 12838 3562
use ota3  X5
timestamp 1729011116
transform 1 0 56242 0 1 9260
box -22 -2458 12838 3562
use ota3  X6
timestamp 1729011116
transform 1 0 69190 0 1 9222
box -22 -2458 12838 3562
use ota3  X7
timestamp 1729011116
transform 0 1 84752 -1 0 12594
box -22 -2458 12838 3562
use ota3  X8
timestamp 1729011116
transform 1 0 69162 0 1 3144
box -22 -2458 12838 3562
use ota3  X9
timestamp 1729011116
transform 1 0 56222 0 1 3126
box -22 -2458 12838 3562
use ota3  X10
timestamp 1729011116
transform 1 0 43254 0 1 3146
box -22 -2458 12838 3562
use ota3  X11
timestamp 1729011116
transform 1 0 30250 0 1 3202
box -22 -2458 12838 3562
use ota3  X12
timestamp 1729011116
transform 1 0 17300 0 1 3258
box -22 -2458 12838 3562
use ota3  X13
timestamp 1729011116
transform 1 0 4352 0 1 3258
box -22 -2458 12838 3562
<< labels >>
flabel via1 16838 -998 17038 -798 0 FreeSans 256 0 0 0 GND
port 3 nsew
flabel via1 4544 -1610 4744 -1410 0 FreeSans 256 0 0 0 VIN
port 11 nsew
flabel metal1 13350 1054 13550 1254 0 FreeSans 256 0 0 0 I0
port 10 nsew
flabel metal1 26302 1056 26502 1256 0 FreeSans 256 0 0 0 I1
port 9 nsew
flabel metal1 39248 998 39448 1198 0 FreeSans 256 0 0 0 I2
port 8 nsew
flabel metal1 52252 946 52452 1146 0 FreeSans 256 0 0 0 I3
port 7 nsew
flabel metal1 65222 922 65422 1122 0 FreeSans 256 0 0 0 I4
port 6 nsew
flabel metal1 78160 940 78360 1140 0 FreeSans 256 0 0 0 I5
port 5 nsew
flabel via1 17510 9822 17710 10022 0 FreeSans 256 0 0 0 C5
port 12 nsew
flabel metal1 30494 9786 30694 9986 0 FreeSans 256 0 0 0 C4
port 13 nsew
flabel via1 43484 9748 43684 9948 0 FreeSans 256 0 0 0 C3
port 14 nsew
flabel metal1 56414 9672 56614 9872 0 FreeSans 256 0 0 0 C2
port 15 nsew
flabel via1 69364 9634 69564 9834 0 FreeSans 256 0 0 0 C1
port 16 nsew
flabel metal1 87000 4598 87200 4798 0 FreeSans 256 0 0 0 VOUT
port 2 nsew
flabel via1 4990 6640 5190 6840 0 FreeSans 256 0 0 0 IOTA
port 1 nsew
flabel via1 6188 12806 6388 13006 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel via1 87228 1398 87428 1598 0 FreeSans 256 0 0 0 VSS
port 4 nsew
<< end >>
