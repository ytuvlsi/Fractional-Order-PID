magic
tech sky130A
magscale 1 2
timestamp 1729526829
<< viali >>
rect 52930 98090 52970 99124
rect 53672 95228 54748 95266
rect 57472 94930 57508 95068
rect 54418 94734 57512 94770
rect 51568 94526 51728 94566
rect 45272 92344 45440 92378
rect 45098 13116 45134 14000
<< metal1 >>
rect 26378 123146 27810 123188
rect 26378 121776 36174 123146
rect 26378 110282 27810 121776
rect 47326 118968 47526 119168
rect 60318 118932 60518 119132
rect 73298 118898 73498 119098
rect 86232 118820 86432 119020
rect 99174 118780 99374 118980
rect 26378 110176 27824 110282
rect 43168 110202 43368 110402
rect 56120 110200 56320 110400
rect 26394 98718 27824 110176
rect 69068 110144 69268 110344
rect 82070 110092 82270 110292
rect 95038 110068 95238 110268
rect 107976 110088 108176 110288
rect 41270 108126 41280 109602
rect 41604 108126 41614 109602
rect 74958 108140 74968 109602
rect 78204 108140 78214 109602
rect 30054 102364 30064 104614
rect 32226 102364 32236 104614
rect 34604 102280 34614 103854
rect 36252 102280 36262 103854
rect 38200 102238 39024 107944
rect 39266 104398 39386 105198
rect 40002 104398 40012 105198
rect 39266 102834 39402 104398
rect 117798 103594 118986 113956
rect 39616 102378 39660 102458
rect 38200 102174 39080 102238
rect 38202 102054 39080 102174
rect 26394 97594 30266 98718
rect 38202 98680 39014 102054
rect 42452 101988 118990 103594
rect 49390 99800 49400 100134
rect 49802 99800 49812 100134
rect 53762 99288 54154 99290
rect 41262 99134 52976 99136
rect 38452 97986 38652 98186
rect 41252 98086 41262 99134
rect 41580 99124 52976 99134
rect 41580 98090 52930 99124
rect 52970 98090 52976 99124
rect 53752 99090 53762 99288
rect 54220 99090 54230 99288
rect 53068 98126 53770 98560
rect 56000 98538 56222 98848
rect 57212 98666 58206 98668
rect 57212 98464 58208 98666
rect 41580 98086 52976 98090
rect 45272 92384 45440 98086
rect 51786 98078 52976 98086
rect 46416 96284 46426 97192
rect 47284 96284 47294 97192
rect 51786 95346 52972 98078
rect 53200 95438 54104 97234
rect 53200 95358 54134 95438
rect 57604 95430 58208 98464
rect 57602 95362 58208 95430
rect 51568 95272 52972 95346
rect 51568 95266 54760 95272
rect 51568 95228 53672 95266
rect 54748 95228 54760 95266
rect 51568 95114 54760 95228
rect 51568 95068 57518 95114
rect 51568 94930 57472 95068
rect 57508 94930 57518 95068
rect 57602 94964 58034 95362
rect 51568 94782 57518 94930
rect 51568 94572 52456 94782
rect 54406 94776 57518 94782
rect 54406 94770 57524 94776
rect 54406 94734 54418 94770
rect 57512 94734 57524 94770
rect 54406 94728 57524 94734
rect 51556 94566 52456 94572
rect 51556 94526 51568 94566
rect 51728 94526 52456 94566
rect 51556 94520 51740 94526
rect 54452 94402 54884 94644
rect 58352 94568 58786 95036
rect 51616 94018 54884 94402
rect 51616 94012 54922 94018
rect 51616 94006 54608 94012
rect 54808 93980 54922 94012
rect 55120 93800 55130 94276
rect 55658 93800 55668 94276
rect 55128 93764 55658 93800
rect 45260 92378 45452 92384
rect 45260 92344 45272 92378
rect 45440 92344 45452 92378
rect 45260 92338 45452 92344
rect 48054 92330 51684 92734
rect 48058 92242 48264 92330
rect 45318 91812 48264 92242
rect 54792 91520 55218 91786
rect 47880 90632 48302 90904
rect 54836 90370 55036 90570
rect 47426 88470 47436 88710
rect 47960 88470 47970 88710
rect 41864 88066 42064 88266
rect 45310 87918 49528 88400
rect 33174 79266 33374 79466
rect 41884 75126 42084 75326
rect 42584 73178 42594 76198
rect 44000 73178 44010 76198
rect 33138 66320 33338 66520
rect 41868 62158 42068 62358
rect 33056 53388 33256 53588
rect 41808 49152 42008 49352
rect 33024 40406 33224 40606
rect 41754 36208 41954 36408
rect 32970 27408 33170 27608
rect 41756 23258 41956 23458
rect 44876 14462 45076 14662
rect 45092 14006 45140 14012
rect 43998 14000 45142 14006
rect 43998 13116 45098 14000
rect 45134 13116 45142 14000
rect 43998 13110 45142 13116
rect 45092 13104 45140 13110
rect 46018 13078 49524 87918
rect 75832 74258 75842 75562
rect 77300 74258 77310 75562
rect 45230 12592 49648 13078
<< via1 >>
rect 41280 108126 41604 109602
rect 74968 108140 78204 109602
rect 30064 102364 32226 104614
rect 34614 102280 36252 103854
rect 39386 104398 40002 105198
rect 49400 99800 49802 100134
rect 41262 98086 41580 99134
rect 53762 99090 54220 99288
rect 46426 96284 47284 97192
rect 55130 93800 55658 94276
rect 47436 88470 47960 88710
rect 42594 73178 44000 76198
rect 75842 74258 77300 75562
<< metal2 >>
rect 30062 115386 35142 116066
rect 30064 104624 32200 115386
rect 41280 109602 41604 109612
rect 74968 109604 78204 109612
rect 74968 109602 78206 109604
rect 78204 108140 78206 109602
rect 74968 108130 78206 108140
rect 41280 108116 41604 108126
rect 39386 105206 40002 105208
rect 39386 105198 49812 105206
rect 26394 104612 28772 104622
rect 30064 104614 32226 104624
rect 25982 102388 26394 104612
rect 28772 102388 30064 104612
rect 26394 102366 28772 102376
rect 32226 102388 32246 104612
rect 40002 104398 49812 105198
rect 39386 104394 49812 104398
rect 39386 104388 40002 104394
rect 34614 103854 36252 103864
rect 30064 102354 32226 102364
rect 39528 102580 39620 102590
rect 39528 102368 39620 102378
rect 34614 102270 36252 102280
rect 41262 99144 41564 100234
rect 48386 100184 49802 104394
rect 48386 100134 53228 100184
rect 48386 99800 49400 100134
rect 49802 99800 53228 100134
rect 48386 99298 53228 99800
rect 48386 99288 54220 99298
rect 41262 99134 41580 99144
rect 48386 99090 53762 99288
rect 48386 99080 54220 99090
rect 48390 99076 54220 99080
rect 48390 99074 53228 99076
rect 41262 98076 41580 98086
rect 46426 97192 47284 97202
rect 46426 96274 47284 96284
rect 51882 94446 53198 99074
rect 54280 99002 54410 99012
rect 54280 98794 54410 98804
rect 51876 94384 53198 94446
rect 51876 94276 55660 94384
rect 51876 93960 55130 94276
rect 47710 89050 47934 89060
rect 47710 88898 47934 88908
rect 47428 88710 47962 88722
rect 47428 88470 47436 88710
rect 47960 88470 47962 88710
rect 47428 88422 47962 88470
rect 51876 88422 52644 93960
rect 55658 93960 55660 94276
rect 55130 93790 55658 93800
rect 55172 93508 55376 93518
rect 55172 93364 55376 93374
rect 74970 92014 78206 108130
rect 74968 92004 78216 92014
rect 74968 91504 78216 91514
rect 47428 87794 52644 88422
rect 51876 87784 52644 87794
rect 36080 84512 36600 84522
rect 36080 81982 36600 81992
rect 42594 76198 44000 76208
rect 48388 76170 49132 76180
rect 44000 73192 48388 76166
rect 74970 76166 78206 91504
rect 49132 75562 78224 76166
rect 49132 74258 75842 75562
rect 77300 74258 78224 75562
rect 49132 73192 78224 74258
rect 44000 73178 78224 73192
rect 42594 73168 44000 73178
rect 74970 73174 78206 73178
<< via2 >>
rect 41280 108126 41604 109602
rect 26394 102376 28772 104612
rect 34614 102280 36252 103854
rect 39528 102378 39620 102580
rect 46426 96284 47284 97192
rect 54280 98804 54410 99002
rect 47710 88908 47934 89050
rect 55172 93374 55376 93508
rect 74968 91514 78216 92004
rect 36080 81992 36600 84512
rect 48388 73192 49132 76170
<< metal3 >>
rect 26384 104612 28782 104617
rect 26384 102376 26394 104612
rect 28772 102376 28782 104612
rect 34372 104004 36394 111250
rect 41270 109602 41614 109607
rect 41270 108126 41280 109602
rect 41604 108126 41614 109602
rect 41270 108121 41614 108126
rect 26384 102371 28782 102376
rect 34362 102190 34372 104004
rect 36418 102190 36428 104004
rect 39428 102328 39438 102656
rect 39726 102328 39736 102656
rect 41276 101890 41602 108121
rect 54212 98732 54222 99012
rect 54422 98732 54432 99012
rect 46416 97192 47294 97197
rect 46416 96284 46426 97192
rect 47284 96284 47294 97192
rect 56602 96862 57202 96864
rect 56016 96496 57202 96862
rect 46416 96279 47294 96284
rect 55120 93364 55130 93692
rect 55418 93364 55428 93692
rect 56602 91984 57202 96496
rect 74958 92004 78226 92009
rect 74958 91984 74968 92004
rect 53572 91540 74968 91984
rect 56602 91538 57202 91540
rect 74958 91514 74968 91540
rect 78216 91514 78226 92004
rect 74958 91509 78226 91514
rect 47672 88858 47682 89062
rect 47948 88858 47958 89062
rect 36070 84512 36610 84517
rect 36070 81992 36080 84512
rect 36600 81992 36610 84512
rect 36070 81987 36610 81992
rect 48388 76175 49134 90880
rect 48378 76170 49142 76175
rect 48378 73192 48388 76170
rect 49132 73192 49142 76170
rect 48378 73187 49142 73192
<< via3 >>
rect 26394 102376 28772 104612
rect 34372 103854 36418 104004
rect 34372 102280 34614 103854
rect 34614 102280 36252 103854
rect 36252 102280 36418 103854
rect 34372 102190 36418 102280
rect 39438 102580 39726 102656
rect 39438 102378 39528 102580
rect 39528 102378 39620 102580
rect 39620 102378 39726 102580
rect 39438 102328 39726 102378
rect 54222 99002 54422 99012
rect 54222 98804 54280 99002
rect 54280 98804 54410 99002
rect 54410 98804 54422 99002
rect 54222 98732 54422 98804
rect 46426 96284 47284 97192
rect 55130 93508 55418 93692
rect 55130 93374 55172 93508
rect 55172 93374 55376 93508
rect 55376 93374 55418 93508
rect 55130 93364 55418 93374
rect 47682 89050 47948 89062
rect 47682 88908 47710 89050
rect 47710 88908 47934 89050
rect 47934 88908 47948 89050
rect 47682 88858 47948 88908
rect 36080 81992 36600 84512
<< metal4 >>
rect 26393 104612 28773 104613
rect 26393 102376 26394 104612
rect 28772 104600 28773 104612
rect 28772 102376 28804 104600
rect 34371 104004 36419 104005
rect 34371 103980 34372 104004
rect 26393 102375 28804 102376
rect 26398 84516 28804 102375
rect 34368 102190 34372 103980
rect 36418 102190 36419 104004
rect 39437 102656 39727 102657
rect 39437 102328 39438 102656
rect 39726 102328 39727 102656
rect 39437 102327 39727 102328
rect 34368 102189 36419 102190
rect 34368 96978 36412 102189
rect 54221 99012 54423 99013
rect 54422 98732 54423 99012
rect 54221 98731 54423 98732
rect 46425 97192 47285 97193
rect 46425 96284 46426 97192
rect 47284 96284 47285 97192
rect 46425 96283 47285 96284
rect 55129 93692 55419 93693
rect 55129 93364 55130 93692
rect 55418 93364 55419 93692
rect 55129 93363 55419 93364
rect 26398 84513 36598 84516
rect 26398 84512 36601 84513
rect 26398 81992 36080 84512
rect 36600 81992 36601 84512
rect 26398 81991 36601 81992
rect 26398 81990 36598 81991
<< via4 >>
rect 39438 102328 39726 102656
rect 54068 98732 54222 99012
rect 54222 98732 54422 99012
rect 46426 96284 47284 97192
rect 55130 93364 55418 93692
rect 47666 89062 47966 89066
rect 47666 88858 47682 89062
rect 47682 88858 47948 89062
rect 47948 88858 47966 89062
rect 47666 88792 47966 88858
<< metal5 >>
rect 39524 102680 47310 102750
rect 39414 102656 47310 102680
rect 39414 102328 39438 102656
rect 39726 102330 47310 102656
rect 39726 102328 39750 102330
rect 39414 102304 39750 102328
rect 46426 99012 47302 102330
rect 54044 99012 54446 99036
rect 46424 98732 54068 99012
rect 54422 98732 54446 99012
rect 46424 98708 54446 98732
rect 46424 98600 54420 98708
rect 46426 97216 47302 98600
rect 46402 97192 47308 97216
rect 46402 96494 46426 97192
rect 46392 96284 46426 96494
rect 47284 96494 47308 97192
rect 47284 96284 47314 96494
rect 46392 93720 47314 96284
rect 46392 93692 55446 93720
rect 46392 93364 55130 93692
rect 55418 93364 55446 93692
rect 46392 93194 55446 93364
rect 47642 89066 48198 93194
rect 47642 88792 47666 89066
rect 47966 88792 48198 89066
rect 47642 88766 48198 88792
use opamp  X1
timestamp 1729086831
transform 1 0 37658 0 1 100478
box 1158 -860 7738 4108
use opamp  X2
timestamp 1729086831
transform 1 0 52410 0 1 96906
box 1158 -860 7738 4108
use opamp  X3
timestamp 1729086831
transform 0 -1 49818 1 0 87042
box 1158 -860 7738 4108
use opamp  X4
timestamp 1729086831
transform 0 1 53276 -1 0 95376
box 1158 -860 7738 4108
use Fractional_diff  X5
timestamp 1729526722
transform 0 -1 43008 1 0 9906
box 3200 -2404 88812 14016
use Fractional_diff  X6
timestamp 1729526722
transform 1 0 29816 0 1 109146
box 3200 -2404 88812 14016
use sky130_fd_pr__res_xhigh_po_0p35_7Z3FVB  XR1
timestamp 1729087846
transform 1 0 53097 0 1 100292
box -201 -2332 201 2332
use sky130_fd_pr__res_xhigh_po_0p35_7Z3FVB  XR2
timestamp 1729087846
transform 0 1 55870 -1 0 95399
box -201 -2332 201 2332
use sky130_fd_pr__res_xhigh_po_0p35_7Z3FVB  XRF
timestamp 1729087846
transform 1 0 45343 0 1 90082
box -201 -2332 201 2332
use sky130_fd_pr__res_xhigh_po_0p35_7Z3FVB  XRW
timestamp 1729087846
transform 0 1 56618 -1 0 94603
box -201 -2332 201 2332
use sky130_fd_pr__res_xhigh_po_0p35_RV8MHK  XRX
timestamp 1729087846
transform 0 1 58193 -1 0 94999
box -201 -757 201 757
use sky130_fd_pr__res_xhigh_po_0p35_JZWPS9  XRY
timestamp 1729087846
transform -1 0 51647 0 -1 93372
box -201 -1230 201 1230
use sky130_fd_pr__res_xhigh_po_0p35_JZWPS9  XRZ
timestamp 1729087846
transform 1 0 45263 0 1 13662
box -201 -1230 201 1230
<< labels >>
flabel metal1 44876 14462 45076 14662 0 FreeSans 256 0 0 0 INPUT
port 6 nsew
flabel metal1 54836 90370 55036 90570 0 FreeSans 256 0 0 0 LOAD
port 7 nsew
flabel metal1 32970 27408 33170 27608 0 FreeSans 256 0 0 0 C5D
port 8 nsew
flabel metal1 33024 40406 33224 40606 0 FreeSans 256 0 0 0 C4D
port 9 nsew
flabel metal1 33056 53388 33256 53588 0 FreeSans 256 0 0 0 C3D
port 10 nsew
flabel metal1 33138 66320 33338 66520 0 FreeSans 256 0 0 0 C2D
port 11 nsew
flabel metal1 33174 79266 33374 79466 0 FreeSans 256 0 0 0 C1D
port 12 nsew
flabel metal1 47326 118968 47526 119168 0 FreeSans 256 0 0 0 C5I
port 13 nsew
flabel metal1 60318 118932 60518 119132 0 FreeSans 256 0 0 0 C4I
port 14 nsew
flabel metal1 73298 118898 73498 119098 0 FreeSans 256 0 0 0 C3I
port 15 nsew
flabel metal1 86232 118820 86432 119020 0 FreeSans 256 0 0 0 C2I
port 16 nsew
flabel metal1 99174 118780 99374 118980 0 FreeSans 256 0 0 0 C1I
port 17 nsew
flabel metal1 38452 97986 38652 98186 0 FreeSans 256 0 0 0 CV
port 31 nsew
flabel metal1 41756 23258 41956 23458 0 FreeSans 256 0 0 0 I0D
port 18 nsew
flabel metal1 41754 36208 41954 36408 0 FreeSans 256 0 0 0 I1D
port 19 nsew
flabel metal1 41808 49152 42008 49352 0 FreeSans 256 0 0 0 I2D
port 20 nsew
flabel metal1 41868 62158 42068 62358 0 FreeSans 256 0 0 0 I3D
port 21 nsew
flabel metal1 41884 75126 42084 75326 0 FreeSans 256 0 0 0 I4D
port 22 nsew
flabel metal1 41864 88066 42064 88266 0 FreeSans 256 0 0 0 I5D
port 23 nsew
flabel metal1 43168 110202 43368 110402 0 FreeSans 256 90 0 0 I0I
port 24 nsew
flabel metal1 56120 110200 56320 110400 0 FreeSans 256 90 0 0 I1I
port 25 nsew
flabel metal1 69068 110144 69268 110344 0 FreeSans 256 90 0 0 I2I
port 26 nsew
flabel metal1 82070 110092 82270 110292 0 FreeSans 256 90 0 0 I3I
port 27 nsew
flabel metal1 95038 110068 95238 110268 0 FreeSans 256 90 0 0 I4I
port 29 nsew
flabel metal1 107976 110088 108176 110288 0 FreeSans 256 90 0 0 I5I
port 30 nsew
flabel via1 31014 103462 31214 103662 0 FreeSans 256 0 0 0 IOTA
port 5 nsew
flabel via1 46752 96694 46952 96894 0 FreeSans 256 0 0 0 IOP
port 4 nsew
flabel via1 76496 74864 76696 75064 0 FreeSans 256 0 0 0 GND
port 3 nsew
flabel via1 49524 99880 49724 100080 0 FreeSans 256 0 0 0 VDD
port 1 nsew
flabel metal1 27030 110904 27230 111104 0 FreeSans 256 0 0 0 VCC
port 0 nsew
flabel via1 35372 103184 35572 103384 0 FreeSans 256 0 0 0 VSS
port 2 nsew
<< end >>
